** sch_path: /home/shaaru/Inv_test.sch
**.subckt Inv_test vout
*.opin vout
x1 vdd vin vout GND inv_vtc
vdd vdd GND 1.8
vin vin GND PULSE(0 1.8 0 .1n .1n 10n 20n 10)
C1 vout GND 10f m=1
**** begin user architecture code

.lib /home/shaaru/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.dc Vin 0 2 1m
.tran .8n 40n
.save all
.end

**** end user architecture code
**.ends

* expanding   symbol:  /home/shaaru/inv_vtc.sym # of pins=4
** sym_path: /home/shaaru/inv_vtc.sym
** sch_path: /home/shaaru/inv_vtc.sch
.subckt inv_vtc vdd vin vout gnd
*.ipin vin
*.ipin vdd
*.ipin gnd
*.opin vout
XM2 vout vin vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 vout vin gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
