* NGSPICE file created from Inv.ext - technology: sky130A
.lib "/home/shaaru/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt"

.subckt Inv in out vdd vss
X0 out in vss vss sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.45 ps=2.9 w=1 l=0.15
X1 out in vdd vdd sky130_fd_pr__pfet_01v8 ad=0.9225 pd=5 as=0.9225 ps=5 w=2.05 l=0.15
.ends Inv

Xinv in out vdd vss Inv

Vdd vdd 0 1.8
Vss vss 0 0

Vin in 0 PULSE(0 1.8 0 1n 1n 10n 20n)

.tran 0.1n 100n

.control
run 
plot v(in) v(out)
.endc

.end
