** sch_path: /home/shaaru/pmos_dc_sweep.sch
**.subckt pmos_dc_sweep
Vgs net2 net1 1.8
Vds net2 GND 0
XM2 GND net1 net2 net2 sky130_fd_pr__pfet_01v8 L=0.15 W=2.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code

.lib /home/shaaru/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.dc Vds 0 2.2 1m
.save all
.end

**** end user architecture code
**.ends
.GLOBAL GND
.end
