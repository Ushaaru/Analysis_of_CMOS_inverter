magic
tech sky130A
timestamp 1715958284
<< nwell >>
rect 0 350 300 770
<< nmos >>
rect 140 200 155 300
<< pmos >>
rect 140 400 155 605
<< ndiff >>
rect 95 290 140 300
rect 95 210 105 290
rect 125 210 140 290
rect 95 200 140 210
rect 155 290 200 300
rect 155 210 170 290
rect 190 210 200 290
rect 155 200 200 210
<< pdiff >>
rect 95 595 140 605
rect 95 410 105 595
rect 125 410 140 595
rect 95 400 140 410
rect 155 595 200 605
rect 155 410 170 595
rect 190 410 200 595
rect 155 400 200 410
<< ndiffc >>
rect 105 210 125 290
rect 170 210 190 290
<< pdiffc >>
rect 105 410 125 595
rect 170 410 190 595
<< psubdiff >>
rect 85 140 210 155
rect 85 110 105 140
rect 190 110 210 140
rect 85 95 210 110
<< nsubdiff >>
rect 65 710 225 720
rect 65 690 80 710
rect 210 690 225 710
rect 65 680 225 690
<< psubdiffcont >>
rect 105 110 190 140
<< nsubdiffcont >>
rect 80 690 210 710
<< poly >>
rect 140 605 155 655
rect 140 375 155 400
rect 100 365 155 375
rect 100 345 110 365
rect 130 345 155 365
rect 100 335 155 345
rect 210 365 250 375
rect 210 345 220 365
rect 240 345 250 365
rect 210 335 250 345
rect 140 300 155 335
rect 140 175 155 200
<< polycont >>
rect 110 345 130 365
rect 220 345 240 365
<< locali >>
rect 65 715 225 720
rect 65 710 125 715
rect 161 710 225 715
rect 65 690 80 710
rect 210 690 225 710
rect 65 685 125 690
rect 161 685 225 690
rect 65 680 225 685
rect 100 605 135 680
rect 95 595 135 605
rect 95 410 105 595
rect 125 410 135 595
rect 95 400 135 410
rect 160 595 200 605
rect 160 410 170 595
rect 190 410 200 595
rect 160 375 200 410
rect 100 365 140 375
rect 100 345 110 365
rect 130 345 140 365
rect 100 335 140 345
rect 160 365 250 375
rect 160 345 220 365
rect 240 345 250 365
rect 160 335 250 345
rect 95 290 135 300
rect 95 210 105 290
rect 125 261 135 290
rect 160 290 200 335
rect 125 210 140 261
rect 95 200 140 210
rect 160 210 170 290
rect 190 210 200 290
rect 160 200 200 210
rect 105 155 140 200
rect 85 145 210 155
rect 85 140 130 145
rect 165 140 210 145
rect 85 110 105 140
rect 190 110 210 140
rect 85 106 130 110
rect 165 106 210 110
rect 85 95 210 106
<< viali >>
rect 125 710 161 715
rect 125 690 161 710
rect 125 685 161 690
rect 110 345 130 365
rect 220 345 240 365
rect 130 140 165 145
rect 130 110 165 140
rect 130 106 165 110
<< metal1 >>
rect -105 715 401 720
rect -105 685 125 715
rect 161 685 401 715
rect -105 679 401 685
rect 20 365 140 375
rect 20 345 110 365
rect 130 345 140 365
rect 20 335 140 345
rect 160 365 400 375
rect 160 345 220 365
rect 240 345 400 365
rect 160 335 400 345
rect -69 156 366 179
rect -71 145 365 156
rect -71 106 130 145
rect 165 106 365 145
rect -71 93 365 106
<< labels >>
rlabel metal1 345 700 345 700 1 vdd
rlabel metal1 305 130 305 130 1 vss
rlabel metal1 375 340 390 365 1 out
rlabel metal1 30 345 45 365 1 in
<< end >>
