** sch_path: /home/shaaru/Dc_sweep.sch
**.subckt Dc_sweep
XM1 Vds Vgs GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vgs Vgs GND 0
Vds Vds GND 0
**** begin user architecture code

.lib /home/shaaru/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.dc Vgs 0 1.8 1m Vds 0 1.8 .5
.save all
.end

**** end user architecture code
**.ends
.GLOBAL GND
.end
